
class hello_world extends uvm_test;
endclass // hello_world
