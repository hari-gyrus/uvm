// ********************************************************************************
// Copyright (c) 2017-2018: Gyrus, Inc
// 
// This file can not be copied and/or distributed without the express permission 
// of Gyrus, Inc. Subject to terms of license agreement - Check "LICENSE" which 
// comes with this distribution for more information.
// ********************************************************************************

class ocp_config;

   // virtual interfaces
   virtual clk_rst_if clk_rst_vif;
   virtual ocp_if     ocp_vif;

endclass // ocp_config

