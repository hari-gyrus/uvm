// ********************************************************************************
// Copyright (c) 2017-2018: Gyrus, Inc
// 
// This file can not be copied and/or distributed without the express permission 
// of Gyrus, Inc. Subject to terms of license agreement - Check "LICENSE" which 
// comes with this distribution for more information.
// ********************************************************************************

//
// ocp_sequencer - ocp slave sequencer
//

typedef uvm_sequencer #(ocp_transaction) ocp_slave_sequencer;

