hari@Haris-MacBook-Pro.local.43377