// ********************************************************************************
// Copyright (c) 2017-2018: Gyrus, Inc
// 
// This file can not be copied and/or distributed without the express permission 
// of Gyrus, Inc. Subject to terms of license agreement - Check "LICENSE" which 
// comes with this distribution for more information.
// ********************************************************************************

package tb_pkg;

  `include "defines.sv"
  `include "ocp_config.sv"
  `include "axi_config.sv"

endpackage // pkg
   
   
