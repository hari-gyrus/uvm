
module design (dut_if d_if);

endmodule // design

